localparam
DECINVALID = 0,
DECREGRS = 1,
DECREGRT = 2,
DECREGFS = 3,
DECREGFT = 4,
DECZIMM = 5,
DECSIMM = 6,
DECALU = 7, /* 5 bit */
DECSETRD = 12,
DECSETRT = 13,
DECMEMRD = 14,
DECMEMWR = 15,
DECSIGNED = 16,
DECSHIMM = 17, /* 2 bit with DECSHIMM32 */
DECSHIMM32 = 18,
DECTARGR = 19, /* 6 bit */
DECLOAD = 25,
DECSZ = 26, /* 4 bit, DECDWORD highest bit */
DECDWORD = 29,
DECLLSC = 30,
DECSTORE = 31,
DECCOND = 32, /* 3 bit */
DECBRANCH = 35,
DECLIKELY = 36,
DECLINK = 37,
DECJUMP = 38,
DECJUMPREG = 39,
DECPANIC = 40,
DECWHY = 41, /* 5 bit */
DECSYSCALL = 46,
DECBREAK = 47,
DECSETFD = 48,
DECSETFT = 49,
DECCACHE = 50,
DECDCACHE = 51,
DECCACHEOP = 52, /* 3 bit */
DECERET = 55,

ALUNOP = 0,
ALUADD = 1,
ALUSUB = 2,
ALUAND = 3,
ALUOR = 4,
ALUNOR = 5,
ALUXOR = 6,
ALUSLL = 7,
ALUSRL = 8,
ALUSRA = 9,
ALUMUL = 10,
ALUDIV = 11,
ALULUI = 12,
ALUADDIMM = 13,
ALUSLT = 14,

CONDAL = 0,
CONDEQ = 1,
CONDNE = 2,
CONDGE = 3,
CONDGT = 4,
CONDLE = 5,
CONDLT = 6,

SZWORD = 0,
SZBYTE = 1,
SZHALF = 2,
SZLEFT = 3,
SZRIGHT = 4,
SZDWORD = 8,
SZDLEFT = 11,
SZDRIGHT = 12,

WHYINTR = 5'h0,
WHYTLBM = 5'h1,
WHYTLBL = 5'h2,
WHYTLBS = 5'h3,
WHYADEL = 5'h4,
WHYADES = 5'h5,
WHYIBE = 5'h6,
WHYDBE = 5'h7,
WHYSYSC = 5'h8,
WHYBRPT = 5'h9,
WHYRSVD = 5'h10,
WHYCPU = 5'h11,
WHYOVFL = 5'h12,
WHYTRAP = 5'h13,
WHYFPE = 5'h15,
WHYWAT = 5'h23,
WHYRST = 5'h31,
WHYNMI = 5'h30,
WHYIADE = 5'h29,
WHYITLB = 5'h28,

/* Status */
IE = 0,
EXL = 1,
ERL = 2,
KSU = 3,
UX = 5,
SX = 6,
KX = 7,
IM = 8,
SR = 20,
TS = 21,
BEV = 22,
RE = 25,
FR = 26,
RP = 27,
CU = 28,

KERN = 0,
SUPR = 1,
USER = 2,

/* CAUSE */
IP = 8,
BD = 31,

/* Config */
K0 = 0,
BE = 15,
EP = 24
;
