`timescale 1 ns / 1 ps
`default_nettype none

`define DECMAX 50
