localparam
DECINVALID = 0,
DECREGRS = 1,
DECREGRT = 2,
DECREGFS = 3,
DECREGFT = 4,
DECZIMM = 5,
DECSIMM = 6,
DECALU = 7, /* 5 bit */
DECSETRD = 12,
DECSETRT = 13,
DECMEMRD = 14,
DECMEMWR = 15,
DECSIGNED = 16,
DECSHIMM = 17, /* 2 bit with DECSHIMM32 */
DECSHIMM32 = 18,
DECTARGR = 19, /* 6 bit */
DECLOAD = 25,
DECSZ = 26, /* 4 bit, DECDWORD highest bit */
DECDWORD = 29,
DECLLSC = 30,
DECSTORE = 31,

ALUNOP = 0,
ALUADD = 1,
ALUSUB = 2,
ALUAND = 3,
ALUOR = 4,
ALUNOR = 5,
ALUXOR = 6,
ALUSLL = 7,
ALUSRL = 8,
ALUSRA = 9,
ALUMUL = 10,
ALUDIV = 11,
ALULUI = 12,
ALUADDIMM = 13,

SZWORD = 0,
SZBYTE = 1,
SZHALF = 2,
SZLEFT = 3,
SZRIGHT = 4,
SZDWORD = 8,
SZDLEFT = 11,
SZDRIGHT = 12,
;
