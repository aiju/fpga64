`include "cpu.vh"

module bus(
	input wire clk,
	input wire bustick,
	
	output wire [31:0] sysadout,
	input wire [4:0] syscmd,
	input wire ereq,
	output wire preq,
	input wire evalid,
	output wire pvalid,
	output wire pmaster,
	input wire eok,
	
	
	
);



endmodule
